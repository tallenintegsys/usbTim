module mem
(
// The $memrd cells have a clock input \CLK, an enable input \EN, an address input \ADDR, and a data output \DATA.
// Clock & reset
input  wire         clk,
input  wire         en,

// PicoRV32 bus interface
input  wire [10:0]  addr,
output reg [7:0]   data);

reg  [7:0] mem[0:1024];

always @(posedge clk) begin
	if (en) begin
		data <= mem[addr];
	end
end

initial begin
	mem[0] = "d";
	mem[1] = "7";
	mem[2] = "b";
	mem[3] = "8";
	mem[4] = "8";
	mem[5] = "c";
	mem[6] = "e";
	mem[7] = "1";
	mem[8] = "6";
	mem[9] = "1";
	mem[10] = "4";
	mem[11] = "3";
	mem[12] = "8";
	mem[13] = "5";
	mem[14] = "5";
	mem[15] = "b";
	mem[16] = "5";
	mem[17] = "a";
	mem[18] = "2";
	mem[19] = "0";
	mem[20] = "d";
	mem[21] = "6";
	mem[22] = "6";
	mem[23] = "a";
	mem[24] = "8";
	mem[25] = "8";
	mem[26] = "a";
	mem[27] = "9";
	mem[28] = "1";
	mem[29] = "f";
	mem[30] = "2";
	mem[31] = "4";
	mem[32] = "b";
	mem[33] = "e";
	mem[34] = "b";
	mem[35] = "0";
	mem[36] = "0";
	mem[37] = "6";
	mem[38] = "f";
	mem[39] = "2";
	mem[40] = "6";
	mem[41] = "d";
	mem[42] = "7";
	mem[43] = "8";
	mem[44] = "1";
	mem[45] = "8";
	mem[46] = "1";
	mem[47] = "2";
	mem[48] = "5";
	mem[49] = "5";
	mem[50] = "e";
	mem[51] = "6";
	mem[52] = "8";
	mem[53] = "4";
	mem[54] = "3";
	mem[55] = "b";
	mem[56] = "e";
	mem[57] = "2";
	mem[58] = "3";
	mem[59] = "b";
	mem[60] = "7";
	mem[61] = "f";
	mem[62] = "b";
	mem[63] = "4";
	mem[64] = "7";
	mem[65] = "0";
	mem[66] = "4";
	mem[67] = "3";
	mem[68] = "2";
	mem[69] = "e";
	mem[70] = "a";
	mem[71] = "7";
	mem[72] = "0";
	mem[73] = "1";
	mem[74] = "3";
	mem[75] = "a";
	mem[76] = "c";
	mem[77] = "2";
	mem[78] = "b";
	mem[79] = "7";
	mem[80] = "c";
	mem[81] = "9";
	mem[82] = "b";
	mem[83] = "5";
	mem[84] = "9";
	mem[85] = "f";
	mem[86] = "e";
	mem[87] = "1";
	mem[88] = "3";
	mem[89] = "a";
	mem[90] = "a";
	mem[91] = "8";
	mem[92] = "1";
	mem[93] = "f";
	mem[94] = "e";
	mem[95] = "2";
	mem[96] = "f";
	mem[97] = "c";
	mem[98] = "6";
	mem[99] = "3";
	mem[100] = "e";
	mem[101] = "f";
	mem[102] = "4";
	mem[103] = "9";
	mem[104] = "e";
	mem[105] = "9";
	mem[106] = "7";
	mem[107] = "6";
	mem[108] = "5";
	mem[109] = "6";
	mem[110] = "b";
	mem[111] = "0";
	mem[112] = "0";
	mem[113] = "c";
	mem[114] = "9";
	mem[115] = "e";
	mem[116] = "3";
	mem[117] = "d";
	mem[118] = "9";
	mem[119] = "f";
	mem[120] = "1";
	mem[121] = "7";
	mem[122] = "e";
	mem[123] = "4";
	mem[124] = "8";
	mem[125] = "3";
	mem[126] = "3";
	mem[127] = "a";
	mem[128] = "e";
	mem[129] = "0";
	mem[130] = "e";
	mem[131] = "8";
	mem[132] = "2";
	mem[133] = "5";
	mem[134] = "a";
	mem[135] = "5";
	mem[136] = "d";
	mem[137] = "4";
	mem[138] = "8";
	mem[139] = "a";
	mem[140] = "5";
	mem[141] = "7";
	mem[142] = "9";
	mem[143] = "a";
	mem[144] = "5";
	mem[145] = "0";
	mem[146] = "c";
	mem[147] = "e";
	mem[148] = "a";
	mem[149] = "2";
	mem[150] = "3";
	mem[151] = "6";
	mem[152] = "7";
	mem[153] = "d";
	mem[154] = "2";
	mem[155] = "4";
	mem[156] = "c";
	mem[157] = "f";
	mem[158] = "d";
	mem[159] = "0";
	mem[160] = "8";
	mem[161] = "e";
	mem[162] = "2";
	mem[163] = "5";
	mem[164] = "6";
	mem[165] = "c";
	mem[166] = "6";
	mem[167] = "e";
	mem[168] = "d";
	mem[169] = "e";
	mem[170] = "9";
	mem[171] = "a";
	mem[172] = "0";
	mem[173] = "c";
	mem[174] = "6";
	mem[175] = "6";
	mem[176] = "7";
	mem[177] = "2";
	mem[178] = "6";
	mem[179] = "7";
	mem[180] = "5";
	mem[181] = "7";
	mem[182] = "6";
	mem[183] = "1";
	mem[184] = "5";
	mem[185] = "1";
	mem[186] = "7";
	mem[187] = "3";
	mem[188] = "e";
	mem[189] = "8";
	mem[190] = "8";
	mem[191] = "2";
	mem[192] = "7";
	mem[193] = "f";
	mem[194] = "6";
	mem[195] = "6";
	mem[196] = "b";
	mem[197] = "1";
	mem[198] = "9";
	mem[199] = "2";
	mem[200] = "3";
	mem[201] = "7";
	mem[202] = "a";
	mem[203] = "b";
	mem[204] = "1";
	mem[205] = "d";
	mem[206] = "5";
	mem[207] = "5";
	mem[208] = "e";
	mem[209] = "3";
	mem[210] = "c";
	mem[211] = "6";
	mem[212] = "6";
	mem[213] = "a";
	mem[214] = "6";
	mem[215] = "b";
	mem[216] = "6";
	mem[217] = "e";
	mem[218] = "0";
	mem[219] = "2";
	mem[220] = "9";
	mem[221] = "3";
	mem[222] = "5";
	mem[223] = "3";
	mem[224] = "a";
	mem[225] = "7";
	mem[226] = "f";
	mem[227] = "2";
	mem[228] = "b";
	mem[229] = "b";
	mem[230] = "1";
	mem[231] = "4";
	mem[232] = "e";
	mem[233] = "2";
	mem[234] = "7";
	mem[235] = "7";
	mem[236] = "7";
	mem[237] = "1";
	mem[238] = "a";
	mem[239] = "6";
	mem[240] = "e";
	mem[241] = "f";
	mem[242] = "a";
	mem[243] = "0";
	mem[244] = "b";
	mem[245] = "8";
	mem[246] = "7";
	mem[247] = "6";
	mem[248] = "8";
	mem[249] = "4";
	mem[250] = "9";
	mem[251] = "f";
	mem[252] = "d";
	mem[253] = "4";
	mem[254] = "5";
	mem[255] = "d";
	mem[256] = "e";
	mem[257] = "e";
	mem[258] = "d";
	mem[259] = "8";
	mem[260] = "1";
	mem[261] = "8";
	mem[262] = "c";
	mem[263] = "6";
	mem[264] = "d";
	mem[265] = "5";
	mem[266] = "e";
	mem[267] = "6";
	mem[268] = "5";
	mem[269] = "3";
	mem[270] = "5";
	mem[271] = "6";
	mem[272] = "f";
	mem[273] = "5";
	mem[274] = "5";
	mem[275] = "9";
	mem[276] = "d";
	mem[277] = "9";
	mem[278] = "4";
	mem[279] = "7";
	mem[280] = "6";
	mem[281] = "8";
	mem[282] = "f";
	mem[283] = "8";
	mem[284] = "e";
	mem[285] = "1";
	mem[286] = "e";
	mem[287] = "8";
	mem[288] = "d";
	mem[289] = "b";
	mem[290] = "c";
	mem[291] = "7";
	mem[292] = "6";
	mem[293] = "c";
	mem[294] = "1";
	mem[295] = "b";
	mem[296] = "7";
	mem[297] = "f";
	mem[298] = "a";
	mem[299] = "1";
	mem[300] = "6";
	mem[301] = "5";
	mem[302] = "6";
	mem[303] = "e";
	mem[304] = "9";
	mem[305] = "5";
	mem[306] = "0";
	mem[307] = "4";
	mem[308] = "c";
	mem[309] = "3";
	mem[310] = "1";
	mem[311] = "b";
	mem[312] = "6";
	mem[313] = "7";
	mem[314] = "d";
	mem[315] = "c";
	mem[316] = "f";
	mem[317] = "8";
	mem[318] = "a";
	mem[319] = "b";
	mem[320] = "1";
	mem[321] = "a";
	mem[322] = "9";
	mem[323] = "4";
	mem[324] = "8";
	mem[325] = "f";
	mem[326] = "3";
	mem[327] = "a";
	mem[328] = "d";
	mem[329] = "6";
	mem[330] = "9";
	mem[331] = "7";
	mem[332] = "1";
	mem[333] = "c";
	mem[334] = "f";
	mem[335] = "3";
	mem[336] = "e";
	mem[337] = "f";
	mem[338] = "f";
	mem[339] = "e";
	mem[340] = "2";
	mem[341] = "4";
	mem[342] = "7";
	mem[343] = "4";
	mem[344] = "0";
	mem[345] = "e";
	mem[346] = "d";
	mem[347] = "1";
	mem[348] = "e";
	mem[349] = "8";
	mem[350] = "3";
	mem[351] = "c";
	mem[352] = "f";
	mem[353] = "4";
	mem[354] = "9";
	mem[355] = "e";
	mem[356] = "6";
	mem[357] = "b";
	mem[358] = "2";
	mem[359] = "e";
	mem[360] = "2";
	mem[361] = "4";
	mem[362] = "7";
	mem[363] = "f";
	mem[364] = "7";
	mem[365] = "6";
	mem[366] = "2";
	mem[367] = "f";
	mem[368] = "e";
	mem[369] = "a";
	mem[370] = "8";
	mem[371] = "3";
	mem[372] = "6";
	mem[373] = "f";
	mem[374] = "c";
	mem[375] = "d";
	mem[376] = "3";
	mem[377] = "2";
	mem[378] = "5";
	mem[379] = "7";
	mem[380] = "3";
	mem[381] = "a";
	mem[382] = "5";
	mem[383] = "f";
	mem[384] = "d";
	mem[385] = "6";
	mem[386] = "8";
	mem[387] = "8";
	mem[388] = "3";
	mem[389] = "d";
	mem[390] = "d";
	mem[391] = "d";
	mem[392] = "d";
	mem[393] = "0";
	mem[394] = "4";
	mem[395] = "2";
	mem[396] = "e";
	mem[397] = "d";
	mem[398] = "8";
	mem[399] = "9";
	mem[400] = "6";
	mem[401] = "8";
	mem[402] = "7";
	mem[403] = "a";
	mem[404] = "d";
	mem[405] = "4";
	mem[406] = "7";
	mem[407] = "c";
	mem[408] = "4";
	mem[409] = "2";
	mem[410] = "7";
	mem[411] = "9";
	mem[412] = "9";
	mem[413] = "1";
	mem[414] = "9";
	mem[415] = "c";
	mem[416] = "9";
	mem[417] = "1";
	mem[418] = "9";
	mem[419] = "3";
	mem[420] = "4";
	mem[421] = "1";
	mem[422] = "0";
	mem[423] = "0";
	mem[424] = "5";
	mem[425] = "e";
	mem[426] = "5";
	mem[427] = "4";
	mem[428] = "6";
	mem[429] = "1";
	mem[430] = "d";
	mem[431] = "e";
	mem[432] = "3";
	mem[433] = "f";
	mem[434] = "9";
	mem[435] = "2";
	mem[436] = "4";
	mem[437] = "6";
	mem[438] = "5";
	mem[439] = "a";
	mem[440] = "e";
	mem[441] = "c";
	mem[442] = "c";
	mem[443] = "1";
	mem[444] = "f";
	mem[445] = "4";
	mem[446] = "8";
	mem[447] = "c";
	mem[448] = "b";
	mem[449] = "5";
	mem[450] = "1";
	mem[451] = "7";
	mem[452] = "a";
	mem[453] = "0";
	mem[454] = "f";
	mem[455] = "1";
	mem[456] = "0";
	mem[457] = "2";
	mem[458] = "1";
	mem[459] = "2";
	mem[460] = "f";
	mem[461] = "e";
	mem[462] = "a";
	mem[463] = "a";
	mem[464] = "6";
	mem[465] = "d";
	mem[466] = "4";
	mem[467] = "1";
	mem[468] = "b";
	mem[469] = "5";
	mem[470] = "1";
	mem[471] = "f";
	mem[472] = "e";
	mem[473] = "b";
	mem[474] = "b";
	mem[475] = "1";
	mem[476] = "1";
	mem[477] = "6";
	mem[478] = "b";
	mem[479] = "e";
	mem[480] = "a";
	mem[481] = "9";
	mem[482] = "0";
	mem[483] = "7";
	mem[484] = "d";
	mem[485] = "b";
	mem[486] = "f";
	mem[487] = "b";
	mem[488] = "0";
	mem[489] = "9";
	mem[490] = "c";
	mem[491] = "6";
	mem[492] = "e";
	mem[493] = "a";
	mem[494] = "c";
	mem[495] = "9";
	mem[496] = "c";
	mem[497] = "a";
	mem[498] = "6";
	mem[499] = "0";
	mem[500] = "7";
	mem[501] = "c";
	mem[502] = "3";
	mem[503] = "f";
	mem[504] = "7";
	mem[505] = "c";
	mem[506] = "4";
	mem[507] = "a";
	mem[508] = "9";
	mem[509] = "2";
	mem[510] = "9";
	mem[511] = "1";
	mem[512] = "a";
	mem[513] = "e";
	mem[514] = "7";
	mem[515] = "a";
	mem[516] = "e";
	mem[517] = "d";
	mem[518] = "d";
	mem[519] = "c";
	mem[520] = "e";
	mem[521] = "b";
	mem[522] = "6";
	mem[523] = "e";
	mem[524] = "3";
	mem[525] = "b";
	mem[526] = "a";
	mem[527] = "2";
	mem[528] = "6";
	mem[529] = "4";
	mem[530] = "9";
	mem[531] = "5";
	mem[532] = "e";
	mem[533] = "7";
	mem[534] = "2";
	mem[535] = "4";
	mem[536] = "d";
	mem[537] = "c";
	mem[538] = "0";
	mem[539] = "0";
	mem[540] = "b";
	mem[541] = "2";
	mem[542] = "2";
	mem[543] = "5";
	mem[544] = "2";
	mem[545] = "f";
	mem[546] = "c";
	mem[547] = "1";
	mem[548] = "b";
	mem[549] = "5";
	mem[550] = "a";
	mem[551] = "1";
	mem[552] = "c";
	mem[553] = "5";
	mem[554] = "8";
	mem[555] = "7";
	mem[556] = "c";
	mem[557] = "4";
	mem[558] = "0";
	mem[559] = "2";
	mem[560] = "5";
	mem[561] = "9";
	mem[562] = "5";
	mem[563] = "1";
	mem[564] = "a";
	mem[565] = "d";
	mem[566] = "7";
	mem[567] = "b";
	mem[568] = "1";
	mem[569] = "0";
	mem[570] = "b";
	mem[571] = "6";
	mem[572] = "b";
	mem[573] = "b";
	mem[574] = "d";
	mem[575] = "c";
	mem[576] = "f";
	mem[577] = "b";
	mem[578] = "b";
	mem[579] = "1";
	mem[580] = "3";
	mem[581] = "d";
	mem[582] = "c";
	mem[583] = "c";
	mem[584] = "7";
	mem[585] = "8";
	mem[586] = "7";
	mem[587] = "1";
	mem[588] = "4";
	mem[589] = "7";
	mem[590] = "8";
	mem[591] = "8";
	mem[592] = "1";
	mem[593] = "d";
	mem[594] = "5";
	mem[595] = "3";
	mem[596] = "e";
	mem[597] = "d";
	mem[598] = "5";
	mem[599] = "5";
	mem[600] = "3";
	mem[601] = "5";
	mem[602] = "8";
	mem[603] = "1";
	mem[604] = "7";
	mem[605] = "3";
	mem[606] = "1";
	mem[607] = "4";
	mem[608] = "5";
	mem[609] = "4";
	mem[610] = "9";
	mem[611] = "4";
	mem[612] = "9";
	mem[613] = "b";
	mem[614] = "1";
	mem[615] = "d";
	mem[616] = "c";
	mem[617] = "1";
	mem[618] = "7";
	mem[619] = "a";
	mem[620] = "b";
	mem[621] = "6";
	mem[622] = "9";
	mem[623] = "8";
	mem[624] = "7";
	mem[625] = "8";
	mem[626] = "6";
	mem[627] = "7";
	mem[628] = "2";
	mem[629] = "5";
	mem[630] = "f";
	mem[631] = "7";
	mem[632] = "d";
	mem[633] = "f";
	mem[634] = "5";
	mem[635] = "d";
	mem[636] = "a";
	mem[637] = "6";
	mem[638] = "b";
	mem[639] = "0";
	mem[640] = "b";
	mem[641] = "8";
	mem[642] = "8";
	mem[643] = "f";
	mem[644] = "e";
	mem[645] = "2";
	mem[646] = "e";
	mem[647] = "4";
	mem[648] = "2";
	mem[649] = "7";
	mem[650] = "5";
	mem[651] = "8";
	mem[652] = "c";
	mem[653] = "b";
	mem[654] = "4";
	mem[655] = "b";
	mem[656] = "f";
	mem[657] = "b";
	mem[658] = "f";
	mem[659] = "c";
	mem[660] = "d";
	mem[661] = "9";
	mem[662] = "a";
	mem[663] = "d";
	mem[664] = "5";
	mem[665] = "1";
	mem[666] = "b";
	mem[667] = "4";
	mem[668] = "d";
	mem[669] = "d";
	mem[670] = "c";
	mem[671] = "9";
	mem[672] = "7";
	mem[673] = "9";
	mem[674] = "5";
	mem[675] = "b";
	mem[676] = "d";
	mem[677] = "1";
	mem[678] = "0";
	mem[679] = "7";
	mem[680] = "9";
	mem[681] = "f";
	mem[682] = "b";
	mem[683] = "c";
	mem[684] = "2";
	mem[685] = "8";
	mem[686] = "c";
	mem[687] = "7";
	mem[688] = "1";
	mem[689] = "d";
	mem[690] = "b";
	mem[691] = "e";
	mem[692] = "c";
	mem[693] = "b";
	mem[694] = "3";
	mem[695] = "7";
	mem[696] = "4";
	mem[697] = "c";
	mem[698] = "d";
	mem[699] = "9";
	mem[700] = "a";
	mem[701] = "7";
	mem[702] = "7";
	mem[703] = "e";
	mem[704] = "6";
	mem[705] = "e";
	mem[706] = "8";
	mem[707] = "e";
	mem[708] = "4";
	mem[709] = "d";
	mem[710] = "1";
	mem[711] = "4";
	mem[712] = "c";
	mem[713] = "a";
	mem[714] = "7";
	mem[715] = "9";
	mem[716] = "0";
	mem[717] = "0";
	mem[718] = "7";
	mem[719] = "3";
	mem[720] = "f";
	mem[721] = "5";
	mem[722] = "d";
	mem[723] = "4";
	mem[724] = "3";
	mem[725] = "7";
	mem[726] = "6";
	mem[727] = "4";
	mem[728] = "d";
	mem[729] = "1";
	mem[730] = "d";
	mem[731] = "9";
	mem[732] = "0";
	mem[733] = "f";
	mem[734] = "e";
	mem[735] = "f";
	mem[736] = "c";
	mem[737] = "3";
	mem[738] = "6";
	mem[739] = "7";
	mem[740] = "3";
	mem[741] = "8";
	mem[742] = "b";
	mem[743] = "c";
	mem[744] = "b";
	mem[745] = "b";
	mem[746] = "f";
	mem[747] = "1";
	mem[748] = "0";
	mem[749] = "9";
	mem[750] = "7";
	mem[751] = "2";
	mem[752] = "b";
	mem[753] = "3";
	mem[754] = "a";
	mem[755] = "3";
	mem[756] = "0";
	mem[757] = "4";
	mem[758] = "f";
	mem[759] = "a";
	mem[760] = "d";
	mem[761] = "5";
	mem[762] = "5";
	mem[763] = "7";
	mem[764] = "7";
	mem[765] = "8";
	mem[766] = "6";
	mem[767] = "4";
	mem[768] = "2";
	mem[769] = "4";
	mem[770] = "a";
	mem[771] = "5";
	mem[772] = "0";
	mem[773] = "5";
	mem[774] = "6";
	mem[775] = "c";
	mem[776] = "1";
	mem[777] = "f";
	mem[778] = "f";
	mem[779] = "5";
	mem[780] = "e";
	mem[781] = "e";
	mem[782] = "1";
	mem[783] = "b";
	mem[784] = "6";
	mem[785] = "2";
	mem[786] = "f";
	mem[787] = "5";
	mem[788] = "f";
	mem[789] = "3";
	mem[790] = "4";
	mem[791] = "5";
	mem[792] = "4";
	mem[793] = "b";
	mem[794] = "b";
	mem[795] = "d";
	mem[796] = "d";
	mem[797] = "5";
	mem[798] = "b";
	mem[799] = "3";
	mem[800] = "2";
	mem[801] = "0";
	mem[802] = "1";
	mem[803] = "2";
	mem[804] = "0";
	mem[805] = "9";
	mem[806] = "b";
	mem[807] = "f";
	mem[808] = "4";
	mem[809] = "6";
	mem[810] = "f";
	mem[811] = "5";
	mem[812] = "b";
	mem[813] = "f";
	mem[814] = "2";
	mem[815] = "f";
	mem[816] = "4";
	mem[817] = "2";
	mem[818] = "f";
	mem[819] = "9";
	mem[820] = "7";
	mem[821] = "e";
	mem[822] = "4";
	mem[823] = "5";
	mem[824] = "6";
	mem[825] = "2";
	mem[826] = "d";
	mem[827] = "7";
	mem[828] = "5";
	mem[829] = "9";
	mem[830] = "e";
	mem[831] = "4";
	mem[832] = "9";
	mem[833] = "a";
	mem[834] = "7";
	mem[835] = "d";
	mem[836] = "4";
	mem[837] = "9";
	mem[838] = "f";
	mem[839] = "e";
	mem[840] = "2";
	mem[841] = "a";
	mem[842] = "3";
	mem[843] = "9";
	mem[844] = "d";
	mem[845] = "e";
	mem[846] = "a";
	mem[847] = "2";
	mem[848] = "e";
	mem[849] = "9";
	mem[850] = "4";
	mem[851] = "d";
	mem[852] = "0";
	mem[853] = "4";
	mem[854] = "3";
	mem[855] = "8";
	mem[856] = "3";
	mem[857] = "b";
	mem[858] = "a";
	mem[859] = "5";
	mem[860] = "b";
	mem[861] = "2";
	mem[862] = "4";
	mem[863] = "e";
	mem[864] = "8";
	mem[865] = "b";
	mem[866] = "5";
	mem[867] = "b";
	mem[868] = "1";
	mem[869] = "9";
	mem[870] = "3";
	mem[871] = "b";
	mem[872] = "4";
	mem[873] = "6";
	mem[874] = "a";
	mem[875] = "1";
	mem[876] = "d";
	mem[877] = "3";
	mem[878] = "1";
	mem[879] = "e";
	mem[880] = "4";
	mem[881] = "1";
	mem[882] = "0";
	mem[883] = "d";
	mem[884] = "a";
	mem[885] = "4";
	mem[886] = "e";
	mem[887] = "5";
	mem[888] = "1";
	mem[889] = "7";
	mem[890] = "b";
	mem[891] = "5";
	mem[892] = "f";
	mem[893] = "3";
	mem[894] = "7";
	mem[895] = "0";
	mem[896] = "9";
	mem[897] = "b";
	mem[898] = "a";
	mem[899] = "0";
	mem[900] = "5";
	mem[901] = "3";
	mem[902] = "7";
	mem[903] = "b";
	mem[904] = "3";
	mem[905] = "6";
	mem[906] = "7";
	mem[907] = "7";
	mem[908] = "b";
	mem[909] = "b";
	mem[910] = "9";
	mem[911] = "9";
	mem[912] = "9";
	mem[913] = "a";
	mem[914] = "9";
	mem[915] = "b";
	mem[916] = "c";
	mem[917] = "7";
	mem[918] = "d";
	mem[919] = "7";
	mem[920] = "b";
	mem[921] = "e";
	mem[922] = "3";
	mem[923] = "d";
	mem[924] = "b";
	mem[925] = "6";
	mem[926] = "4";
	mem[927] = "5";
	mem[928] = "9";
	mem[929] = "4";
	mem[930] = "3";
	mem[931] = "1";
	mem[932] = "0";
	mem[933] = "d";
	mem[934] = "a";
	mem[935] = "1";
	mem[936] = "2";
	mem[937] = "2";
	mem[938] = "b";
	mem[939] = "c";
	mem[940] = "a";
	mem[941] = "9";
	mem[942] = "0";
	mem[943] = "6";
	mem[944] = "6";
	mem[945] = "6";
	mem[946] = "f";
	mem[947] = "6";
	mem[948] = "0";
	mem[949] = "0";
	mem[950] = "0";
	mem[951] = "5";
	mem[952] = "5";
	mem[953] = "9";
	mem[954] = "0";
	mem[955] = "5";
	mem[956] = "7";
	mem[957] = "d";
	mem[958] = "2";
	mem[959] = "1";
	mem[960] = "9";
	mem[961] = "d";
	mem[962] = "c";
	mem[963] = "0";
	mem[964] = "8";
	mem[965] = "f";
	mem[966] = "b";
	mem[967] = "d";
	mem[968] = "3";
	mem[969] = "4";
	mem[970] = "f";
	mem[971] = "2";
	mem[972] = "a";
	mem[973] = "0";
	mem[974] = "6";
	mem[975] = "a";
	mem[976] = "7";
	mem[977] = "3";
	mem[978] = "c";
	mem[979] = "9";
	mem[980] = "c";
	mem[981] = "f";
	mem[982] = "7";
	mem[983] = "0";
	mem[984] = "2";
	mem[985] = "d";
	mem[986] = "5";
	mem[987] = "e";
	mem[988] = "d";
	mem[989] = "d";
	mem[990] = "0";
	mem[991] = "b";
	mem[992] = "1";
	mem[993] = "a";
	mem[994] = "2";
	mem[995] = "2";
	mem[996] = "d";
	mem[997] = "f";
	mem[998] = "0";
	mem[999] = "2";
	mem[1000] = "8";
	mem[1001] = "a";
	mem[1002] = "e";
	mem[1003] = "0";
	mem[1004] = "2";
	mem[1005] = "9";
	mem[1006] = "8";
	mem[1007] = "a";
	mem[1008] = "d";
	mem[1009] = "e";
	mem[1010] = "e";
	mem[1011] = "8";
	mem[1012] = "8";
	mem[1013] = "2";
	mem[1014] = "8";
	mem[1015] = "9";
	mem[1016] = "7";
	mem[1017] = "f";
	mem[1018] = "e";
	mem[1019] = "8";
	mem[1020] = "8";
	mem[1021] = "7";
	mem[1022] = "f";
	mem[1023] = "c";
end
endmodule
